module and_gate(out, a, b);
    output out1;
    input a,b;

    and a1 (out, a, b);
endmodule